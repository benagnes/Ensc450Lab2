.alter xor_x1_a_fall_2
Xxor_x1_a_fall  a_fall   gnd   z    vdd vdds gnd gnds xr    ds=1
.param Cload=2fF

.alter xor_x1_a_fall_10
.param Cload=10fF



.alter xor_x4_a_fall_2
Xxor_x4_a_fall  a_fall   gnd   z    vdd vdds gnd gnds xr    ds=4
.param Cload=2fF

.alter xor_x4_a_fall_10
.param Cload=10fF





.alter xor_x1_b_fall_2
Xxor_x1_b_fall  gnd   a_fall   z    vdd vdds gnd gnds xr    ds=1
.param Cload=2fF

.alter xor_x1_b_fall_10
.param Cload=10fF



.alter xor_x4_b_fall_2
Xxor_x4_b_fall  gnd   a_fall   z    vdd vdds gnd gnds xr    ds=4
.param Cload=2fF

.alter xor_x4_b_fall_10
.param Cload=10fF



.end
