.alter xorlay_x1_a_fall_2
Xxorlay_x1_a_fall  a_fall   gnd   z    vdd vdds gnd gnds xrlay    ds=1
.param Cload=2fF

.alter xorlay_x1_a_fall_10
.param Cload=10fF



.alter xorlay_x4_a_fall_2
Xxorlay_x4_a_fall  a_fall   gnd   z    vdd vdds gnd gnds xrlay    ds=4
.param Cload=2fF

.alter xorlay_x4_a_fall_10
.param Cload=10fF





.alter xorlay_x1_b_fall_2
Xxorlay_x1_b_fall  gnd   a_fall   z    vdd vdds gnd gnds xrlay    ds=1
.param Cload=2fF

.alter xorlay_x1_b_fall_10
.param Cload=10fF



.alter xorlay_x4_b_fall_2
Xxorlay_x4_b_fall  gnd   a_fall   z    vdd vdds gnd gnds xrlay    ds=4
.param Cload=2fF

.alter xorlay_x4_b_fall_10
.param Cload=10fF



.end
